module days

fn test_day_three() {
	run_tests(day_three, [
		TestFixture{read_input(day: 3), '4361', '467835'},
	])
}
