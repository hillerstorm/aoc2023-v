module days

fn test_day_two() {
	run_tests(day_two, [
		TestFixture{read_input(day: 2), '8', '2286'},
	])
}
