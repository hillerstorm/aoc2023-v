module days

fn test_day_five() {
	run_tests(day_five, [
		TestFixture{read_input(day: 5), '35', '46'},
	])
}
