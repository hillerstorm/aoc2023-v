module days

fn test_day_four() {
	run_tests(day_four, [
		TestFixture{read_input(day: 4), '13', '30'},
	])
}
