module days

fn test_day_six() {
	run_tests(day_six, [
		TestFixture{read_input(day: 6), '288', '71503'},
	])
}
